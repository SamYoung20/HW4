//Deliverable 2
module register
  (
  output reg	q,
  input		d,
  input		wrenable,
  input		clk
  );

      always @(posedge clk) begin
          if(wrenable) begin
              q <= d;
          end
      end

endmodule
